module XOR(input logic[2:0] a,b , output logic[2:0] f);
    assign f = a^b;
endmodule