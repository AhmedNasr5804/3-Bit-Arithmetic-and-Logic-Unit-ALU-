module AND(input logic[2:0] a, b, output reg[2:0] y);
    assign y = a & b;
endmodule