module cmp( input logic [2:0] A, output logic [2:0] F);
    assign F = ~A;
endmodule
